package counter_types;

typedef enum logic[1:0] {
  NONE, INC, LOAD
} cmd_t /* verilator public */;

endpackage
