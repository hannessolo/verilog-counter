package alu_types;

typedef enum logic[1:0] {
  ADD,
  SUB,
  OR,
  AND
} alu_t;

endpackage
