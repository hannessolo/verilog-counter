package microaddr;

typedef enum logic[1:0] {
  NONE, INC, LOAD
} cmd /* verilator public */;

endpackage
